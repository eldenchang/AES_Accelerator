PK  ��L               word/numbering.xml��MN�0�O�"��$ 5�
6����X�=��I��q��R$��U��������Kɠ�h��ˈ\3Ȅ.R���x"�uTgT��)9rK���u��J�9�}�Gh�(���9���e%W�.�p�9���/��Ce��N�����tHI�:�%��ܝ$	�`���
���Jv�*ŵ;;�ȥ��-��=Mͥ�b�C�Q+��k��i��dk� f�qk��][�q4a�'Ġ���OϾE�0�t\����vF�ga�F�қ�#���.�y^ꍘ��+�W�
�@�A����rA;���aΊIq�"e�H�R{����U\�Kj�H+�G{E����9��?�X��p�PKICh  =  PK  ��L               word/settings.xml���n�0ǟ`����I6uzX���= #ɶ}A����'ǖդ@�f�H�?�M?>�|q��2%K��R��+�d]�?�?����:����Dgj����cWX���O���D�s�H�*�����+e85u"�[��Jhp��8s�$O�-1�D��ňX
����r}H���a:��3'��p+�t�����נ�m���&�yc ���$x����l�@�-���S�h�0�֫σq"f���)bN	�9C%��0�p܀��+�{l�$���9����`���Ww��m�f�����\k����0. �=��� O03�g���0��8��S�l�ތ˾M#��?�O�Z�}}���m>�`�W ��ܽ�a�^t�	��S���a���~ؘ�/[#� ��s�_���5l~q}��*'7�>����C�C�����qY�w�F�B�\u>��-l�`����Q˃���!hQ[m�M�6Q�m�k�YSÙ<�6�c�W�s�Q�+��Ic?�Wj�PK����  �  PK  ��L               word/fontTable.xml��MN�0�O�"�ۤ��Tv��I��k�4���4?P$��U�������7ZE;AN���j��H��4U��^�,rL
���^8��/�mZ��.
r�R�3V{o�8v���0�X"i�ᕪXm��-x�.����2InX���5d��В:,�A�bYJ.�G��)�G��F�c*���Һ����B��!��6�Ӫ_��)nA�B��Q�TXB.�_�Ł�J&��SZ���w�A�sH�	h�^�nh_�q#�,���ȱ�,�	h���1��z+'���T��!�s��=@�!(�[Q܃��梚�R!�"�cH�Y'�JN��R�#��퉰�cܯ�о����� �= �M��;��X����b�?PK��m y  Z  PK  ��L               word/styles.xmlՖ�n�0��`���MHCQiU��6�ꦵ���c�UǶlʮ~�7$�J� ���~�:���[LGk,�ln�/k��!a������bf���ϭ-V�����M���b52�L1�[��"�m�"���3ӹ�2m�re� _q�x,@��Dom�q�V!��V"YPH\�I��R�)_.	��O�!���S�9Jb�tVі��9p�""T�U3�Q)�~o똖�6�O�P��lFL�B.C!9�J��}�Y)�� S�*���k�3���J&�FC��}ij�2�z!5E�L$�z$	r۞๛/H/7L�Nde�!(�K:D�r��;`k���zٹ�XI�k�����i��9�k��qj�$ODmw���	O>&����rt���P�Ҧ�%�f��~8�j�	@!B�֭$`�o�v��UvB�-S�x;�RMx核n�S��*c��1���ݜ�h�2M�d�����:��� $������[\�{�H�0�d�/��Y׏pn=�~����*�3�q���kg�my���_�H/�l��G��E|ǐ^�m�(���-Z���OV��M~�]�bs^1O;C
�4�h6H5��^�RcsS�]'����o��;��{[ٸ��ﴽ��v|6�{��ɰyӾ����<�^��cGb�b�΍q�O�Jq�e�=/������'��x��x�υם�Ż�s�}Z8���	pN�|2��)q����9=�s���$��}!ڼU���虹N��~�>�t���9Y�N^UǙ�y� f'|��L�u�u���x���w����?PK��E  �  PK  ��L               word/document.xml��n�0ǟ`ڤ�`B���նlӤm���jڅX۲M���gbC���Ҭ�X.
�����;>����۲�XH������a����l���x2�=�MQ�(��+,���gK���*1U�V����ϕ�0d���S�1Օs&J���Ȃ�_?IXɑ"3R�
�0�V�M�JPh%NJ�&�\�M ��I��i!���4�Z��=�FeN�l��C�teވ,Ģ,���|��R��GY���L�\�K�K���U��%�����gcI�me��#��}���N[Km��,�1�T}!3���� n��d�(���[�J�y�D�#�����%�p��j�9��
�;J)A�@�&H�Ȃ�N�\��Z�wj���&��CԶf �?M j�u
��tU���:��W?�?�Mqq���~���QU�j.�N!�!G}N�J�F\���0��Pq�Q��e�6��zq)�1h�����vͱ��*v�
ښ�#Jm��\`����%K�{�.�s2W/�ʴ3:�Zp����ϺS�A���{	��%���!j&�]���4X�j;4t��4z�I����3��H?�3ZG�:�A�C{�SM{�$�~����p4�X̹�P��2����B1�NBv
J�(�P̹�PFNCq�Uc�]��`0� D6��������2�Q�.�����SX�}7�"��I(�;�$-� r��i(N��Ӯz�G0� l��Ǝ�����2�a�.�`'��#}� 39�e��6Nb����v����bf��L��6p�UG�N���{pܬ � M*��0 웵1�9�U��1`@ؙ�\��nm���͊��1'���+��������UG����|���L�8Q�9Ϯk�|��(^���Q�!��+��1cJ�RW��.����s��$˷.s�R,Z��[Uެ8�UR!Q�i�Ԙ4����� PK��.��  A,  PK  ��L               word/_rels/document.xml.rels��Mj�0�O�;��ײ�J��Md[�(���Z#!MJ}���$Ӆ��y�֛͌;�o�w���rH��=�
>����Țj=8B#Fؔ�4����>�BQA��ߥ��C�c�<Rzi\������|��*�_e�f@y�)��������?ٮiz�[g��ﴐ�j1��"+8�?��R���%"2���+�ٙCxZ�qĕ>�U\�9��%!�h��W��5��1xpz��>��7���PK� ���   ,  PK  ��L               _rels/.rels��;�0�p��;Mˀj�!uE� Q��CIx��d` ��h��g��v&7��xǠ�j �W�i���IY8%f���	:�jO8�\v�dB"q���s�S��V��te2�hE.e�4y馮�4��?L�+�W�a	�����H<xy���_�"��13����z����-�x�?PK-h�"�   *  PK  ��L               word/theme/theme1.xml�YKo�6��w toe�V�u�رۭM$n�i���P�@�I|��úa��m�a[�إ�4�:lЯ���)�ΣM��6I���I��È�}"$�q�r.�,Db��4���A�B�BR��ǌǤmM������e��B��\�m+T*Y�m��2�yBbx6�"�
�"�}��o��z��bG���qlo�F�#h���֧�{�b%���]/��SdX�I�Dv�@���-���9TbX*xжj�ǲ�/�%SKh5�~�)�
��щ`X:���͒=翈��zݞS�� ���Rg�췜Δ�ʇ���5�֬�5���j��qW+���\��j+͍zߜ��E�;��J���+���Օf��BF�t�22%d��5#���4f([ˮ�>V�r-���� .V4Fj��� �ŌM�5��'��'�RYHz�&�m}�`����_>{���?=���уG�6P]�q�S�����}��z�݋�_��R����g�����t�������o>�����C>���&9@;<��P��bb�Slā�1Ni�
+�̰�!U��L���{�wC1V� �F��ÅѦ�,��80c���Ivw.��q�LM,�!���� �8 1Q(}��1�ݥ���-�	.�H��u05�d@��Lt�F��IA�w�7[wP�3�M�_EBU`fbIXōW�X�Ȩ1�����UhRrw"��å�H�q��&�[bRQ�:�sط�$�"��{&�̹���{�G�Qg�:�#�)��6WF%x�B�9��K�}�u�ھM�М 铱0���z��&q��+�:��q�;���ϻqC�|���Q�� '�jf�Q/�ͷ�.>}���&��
�}s~ߜ��漬�Ͽ%Ϻ���36��S��2��&�ܐY��`�߇�l����$�a!����Hp�	U�n��dY�$J������wv?�`s��N/���j���rC�l�l�Y uA���i�5.��0'�R�㚥��J�5oB� ��JpV�hH̈��=g0��S�bb��5����{&%��ɵ'ۋ������U��Z��I��i	�Q�d�i0�����kq��UsV95w����j�0��M_��3��n3���`h&�Ӣ�r�C-��Вшxj��lZ<�cE�n��!�z7���N_�N�v�H�j��1�ʦ�̒���b�óq�C6�Գ�����4����5%�\8�6������(�ѶŅ
9t�$�^_������E�b��TW�?�[9����ڡ:�
!۪��fN]����>S�+��wH�	�ջ��o�p�M
Gd���٦������|��g&�y�ͯ�5}m+X}=N�k��f���ҝg~�M����/h�Txlv<��>*�y�x�U�_�8�[�q)���Z��<;j�n,q���^�ٮ����K���!�l�(>��7�z3f��L`��Ef���b�d�rGL[:�w�Q�p�9������N. ��$l�LX�g�HI\?������J��gb�f�s|�E��b���ʛ]f��Ӻ��z����]Vx�6%9Tw�]A�ڳ�]�PK!Z��,  �  PK  ��L               [Content_Types].xml��Mn�0�O�;D�V��EUU�Y�]����O����;	�����e�ͼ�y$O�;�-f�1TjR�U���چU�>��UC��ŀ��#���f��'�B�Uj͜�&�FTƄA�&f,Ǽ�	��Pߍ�����xĭ��M�������p�ZW
Rr� �3U��D<`�g���m��`FG�2��jhmݞ�Jm»L&�������xi)�c�S��d�ޕ�̲;�~@�7�b��J}R��#�A��k �6h|#^X:�L�˃B��_b��e�^�W<�p�/�G��ze��tX'�H����PK3��,  -  PK   ��LICh  =                   word/numbering.xmlPK   ��L����  �               �  word/settings.xmlPK   ��L��m y  Z               �  word/fontTable.xmlPK   ��L��E  �               �  word/styles.xmlPK   ��L��.��  A,               �  word/document.xmlPK   ��L� ���   ,               �  word/_rels/document.xml.relsPK   ��L-h�"�   *               ,  _rels/.relsPK   ��L!Z��,  �                 word/theme/theme1.xmlPK   ��L3��,  -               �  [Content_Types].xmlPK    	 	 B  �    